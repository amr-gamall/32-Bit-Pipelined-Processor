`include "Instruction-Memory/instruction_memory.v"
`include "Data-Memory/Data_Memory.v"
`include "ALU/alu.v"
`include "Register-File/Register-File.v"
`include "Program-Counter/Program_Counter.v"

module dataPath(
    input         rst, clk,

);


endmodule
